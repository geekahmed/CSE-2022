$date
  Sat Nov 21 23:38:34 2020
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module task1tb $end
$var reg 1 ! a $end
$var reg 1 " b $end
$var reg 1 # c $end
$var reg 1 $ d $end
$var reg 1 % e $end
$var reg 1 & f $end
$var reg 1 ' g $end
$var reg 1 ( h $end
$var reg 1 ) i $end
$scope module tree $end
$var reg 1 * a $end
$var reg 1 + b $end
$var reg 1 , c $end
$var reg 1 - d $end
$var reg 1 . e $end
$var reg 1 / f $end
$var reg 1 0 g $end
$var reg 1 1 h $end
$var reg 1 2 i $end
$var reg 1 3 sig1 $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
X!
X"
X#
X$
X%
X&
X'
X(
X)
X*
X+
X,
X-
X.
X/
X0
X1
X2
X3
#1000000
1!
0"
0#
0$
0%
0&
0'
1(
0)
1*
0+
0,
0-
0.
0/
00
11
02
03
#2000000
0!
1"
0(
0*
1+
01
#3000000
0"
1#
0+
1,
#4000000
0#
1$
0,
1-
#5000000
0$
1%
0-
1.
#6000000
0%
1&
0.
1/
#7000000
#8000000
